// Created by Jeevaka Dassanayake on 5/24/18.
//   Copyright (c) 2018 Jeevaka Dassanayake.

`timescale 1ns / 1ps

module BoardTest( input wire clk, input wire [4:0] bt, input wire [7:0] dp, output wire [7:0] ss, output wire [2:0] en );


endmodule
