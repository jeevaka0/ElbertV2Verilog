// Created by Jeevaka Dassanayake on 5/08/18.
//   Copyright (c) 2018 Jeevaka Dassanayake.

`timescale 1ns / 1ps

module DualPriority( input wire [12:1] r, output reg [3:0] first , output reg [3:0] second );

always @*
begin
	casez (r)
		12'b1???????????: first = 4'b1100;
		12'b01??????????: first = 4'b1011;
		12'b001?????????: first = 4'b1010;
		12'b0001????????: first = 4'b1001;
		12'b00001???????: first = 4'b1000;
		12'b000001??????: first = 4'b0111;
		12'b0000001?????: first = 4'b0110;
		12'b00000001????: first = 4'b0101;
		12'b000000001???: first = 4'b0100;
		12'b0000000001??: first = 4'b0011;
		12'b00000000001?: first = 4'b0010;
		12'b000000000001: first = 4'b0001;
		12'b000000000000: first = 4'b0000;
	endcase
end

always @*
begin
	casez (r)
		12'b11??????????: second = 4'b1011;
		12'b101?????????, 12'b011?????????: second = 4'b1010;
		12'b1001????????, 12'b0101????????, 12'b0011????????: second = 4'b1001;
		12'b10001???????, 12'b01001???????, 12'b00101???????, 12'b00011??????? : second = 4'b1000;
		12'b100001??????, 12'b010001??????, 12'b001001??????, 12'b000101??????, 12'b000011?????? : second = 4'b0111;
		12'b1000001?????, 12'b0100001?????, 12'b0010001?????, 12'b0001001?????, 12'b0000101?????, 12'b0000011?????
			: second = 4'b0110;
		12'b10000001????, 12'b01000001????, 12'b00100001????, 12'b00010001????, 12'b00001001????, 12'b00000101????
			, 12'b00000011???? : second = 4'b0101;
		12'b100000001???, 12'b010000001???, 12'b001000001???, 12'b000100001???, 12'b000010001???, 12'b000001001???
			, 12'b000000101???, 12'b000000011??? : second = 4'b0100;
		12'b1000000001??, 12'b0100000001??, 12'b0010000001??, 12'b0001000001??, 12'b0000100001??, 12'b0000010001??
			, 12'b0000001001??, 12'b0000000101??, 12'b0000000011?? : second = 4'b0011;
		12'b10000000001?, 12'b01000000001?, 12'b00100000001?, 12'b00010000001?, 12'b00001000001?, 12'b00000100001?
			, 12'b00000010001?, 12'b00000001001?, 12'b00000000101?, 12'b00000000011? : second = 4'b0010;
		12'b100000000001, 12'b010000000001, 12'b001000000001, 12'b000100000001, 12'b000010000001, 12'b000001000001
			, 12'b000000100001, 12'b000000010001, 12'b000000001001, 12'b000000000101, 12'b000000000011 : second = 4'b0001;
		12'b000000000000, 12'b000000000001, 12'b000000000010, 12'b000000000100, 12'b000000001000, 12'b000000010000
			, 12'b000000100000, 12'b000001000000, 12'b000010000000, 12'b000100000000, 12'b001000000000
			, 12'b010000000000, 12'b100000000000: second = 4'b0000;
	endcase
end

endmodule
